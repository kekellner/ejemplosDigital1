module tabla01POS();


endmodule